module pianocontroller();

endmodule 