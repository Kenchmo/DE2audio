module pianocontroller();












end module 